library verilog;
use verilog.vl_types.all;
entity wrapper_test is
end wrapper_test;
