library verilog;
use verilog.vl_types.all;
entity design_test is
end design_test;
